// imm_generator.v

module imm_generator #(
  parameter DATA_WIDTH = 32
)(
  input [31:0] instruction,

  output reg [DATA_WIDTH-1:0] sextimm
);

wire [6:0] opcode;
assign opcode = instruction[6:0];

always @(*) begin
  case (opcode)
    //////////////////////////////////////////////////////////////////////////
    // TODO : Generate sextimm using instruction (DONE)
    //////////////////////////////////////////////////////////////////////////
    6'b0010011: sextimm = $signed(instruction[31:20]);
    
    default:    sextimm = 32'h0000_0000;
  endcase
end


endmodule
