module branch_control
(
  // current pc
  input branch,
  input check,

  output reg taken 
);

///////////////////////////////////////////////////////////////////////////////
// TODO : You need to do something! (DONE)
//////////////////////////////////////////////////////////////////////////////

always @(*) begin
  taken = branch & check ?  1'b1 : 1'b0;
end

endmodule
